module Prob002_m2014_q4i_spec(output [0:0] out);
    assign out = 1'b0; // always drive logic low
endmodule

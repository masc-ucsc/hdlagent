module Prob003_step_one_spec(output [0:0] one);
    assign one = 1'b1; // Always drive the output 'one' to logic high (1)
endmodule

module Prob007_wire_spec(input [0:0] in, output [0:0] out);
    assign out = in; // Wire behavior: output directly connected to input
endmodule

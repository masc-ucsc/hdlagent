module hex_literal_demo_spec(output [15:0] o);
  assign o = 16'hA55A; // Set output to hexadecimal literal 0xA55A
endmodule

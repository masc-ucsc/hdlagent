module hex_literal_demo (
    output reg [15:0] o
);

assign o = 16'hA55A;

endmodule
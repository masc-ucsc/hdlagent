module priority_encoder
  (
  input [24:0] significand, 
  input [7:0] exp_a, 
  output reg [24:0] Significand, 
  output reg [7:0] exp_sub
  );

// Here insert your combinational logic for the priority encoder

endmodule
module Prob001_zero_spec(output [0:0] zero);
    // Assign constant LOW to the zero output
    assign zero = 1'b0;
endmodule

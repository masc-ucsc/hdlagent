module TopModule(
    input [0:0] in, 
    output [0:0] out
);

assign out = in; // Combinational assignment

endmodule
